package IKA9958_mnemonics;

localparam T1 = 5'b00001;
localparam T2 = 5'b01001;

endpackage : IKA9958_mnemonics
