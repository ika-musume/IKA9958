package IKA9958_mnemonics;

localparam T1 = 5'b00001;
localparam T2 = 5'b01001;
localparam MC = 5'b00010;
localparam G1 = 5'b00000;
localparam G2 = 5'b00100;
localparam G3 = 5'b01000;
localparam G4 = 5'b01100;
localparam G5 = 5'b10000;
localparam G6 = 5'b10100;
localparam G7 = 5'b11100;


endpackage : IKA9958_mnemonics
