module IKA9958_rcc #(parameter CM = 1) (

);

/*
    IKA9958 Reset and Clock Control
*/


endmodule