/*
    IKA9958 Buses

    Lists all interface modules for internal tri-state buses
*/