module IKA9958_st (

);

/*
    IKA9958 Screen Timing
    This module generates all video timing signals
*/








endmodule